----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:11:34 12/28/2016 
-- Design Name: 
-- Module Name:    pc - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pc is

    Port ( a : in  STD_LOGIC_VECTOR (31 downto 0);
           clk : in  STD_LOGIC;
           b : out  STD_LOGIC_VECTOR (31 downto 0));

end pc;

architecture Behavioral of pc is

begin

process (clk,a )

begin 

if rising_edge (clk) 
    then b <= a;

end if ;

end process;
end Behavioral;

